
-- Based on Xilinx Parity Checker Mealy State Machine Example
-- https://www.xilinx.com/support/documentation/university/Vivado-Teaching/HDL-Design/2015x/VHDL/docs-pdf/lab10.pdf
-- Page 10-1 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity separate_state_and_comb_next is
  port (
    iClk                : in std_logic;
    iReset              : in std_logic;
    iData               : in std_logic;
    oParity             : out std_logic :='0'
  ) ;
end entity ; -- separate_state_and_comb_next

architecture rtl of separate_state_and_comb_next is

  type state_type is (S0, S1);
  signal state, next_state : state_type;

  signal parity_comb : std_logic := '0';

begin

  RESET_PROC : process (iClk)
  begin
    if rising_edge(iClk) then
      if (iReset = '1') then
        state <= S0;
      else
        state <= next_state;
      end if;
    end if;
  end process;

  -- Register output without reset
  SYNC_PROC : process (iClk)
  begin
    if rising_edge(iClk) then
      oParity <= parity_comb;
    end if;
  end process;

  NEXT_STATE_DECODE : process (state, iData)
  begin
    parity_comb <= '0';
    case (state) is
      when S0 =>
        if (iData = '1') then
          parity_comb <= '1';
          next_state  <= S1;
        else
          next_state  <= S0;
        end if;
      when S1 =>
        if (iData = '1') then
          next_state  <= S0;
        else
          parity_comb <= '1';
          next_state  <= S1;
        end if;
      when others =>
        next_state <= S0;
    end case;
  end process;

end architecture ; -- rtl
